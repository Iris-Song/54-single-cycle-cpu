`timescale 1ns / 1ps

module clz(
   input  [31:0]clz_in,
   output [31:0]clz_out
    );
    
     assign clz_out = clz_in[31]==1? 32'h00000000:clz_in[30]==1? 32'h00000001:clz_in[29]==1? 32'h00000002:clz_in[28]==1? 32'h00000003:clz_in[27]==1? 32'h00000004:
                      clz_in[26]==1? 32'h00000005:clz_in[25]==1? 32'h00000006:clz_in[24]==1? 32'h00000007:clz_in[23]==1? 32'h00000008:clz_in[22]==1? 32'h00000009:
                      clz_in[21]==1? 32'h0000000a:clz_in[20]==1? 32'h0000000b:clz_in[19]==1? 32'h0000000c:clz_in[18]==1? 32'h0000000d:clz_in[17]==1? 32'h0000000e:
                      clz_in[16]==1? 32'h0000000f:clz_in[15]==1? 32'h00000010:clz_in[14]==1? 32'h00000011:clz_in[13]==1? 32'h00000012:clz_in[12]==1? 32'h00000013:
                      clz_in[11]==1? 32'h00000014:clz_in[10]==1? 32'h00000015:clz_in[9]==1? 32'h00000016:clz_in[8]==1? 32'h00000017:clz_in[7]==1? 32'h00000018:
                      clz_in[6]==1? 32'h00000019:clz_in[5]==1? 32'h0000001a:clz_in[4]==1? 32'h0000001b:clz_in[3]==1? 32'h0000001c:clz_in[2]==1? 32'h0000001d:
                      clz_in[1]==1? 32'h0000001e:clz_in[0]==1? 32'h0000001f:32'h00000020;
     
endmodule
